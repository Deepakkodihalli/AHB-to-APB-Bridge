package pkg;

import uvm_pkg::*;

`include "uvm_macros.svh"

`include "ahb_config.sv"
`include "ahb_trans.sv"
`include "ahb_seqs.sv"
`include "ahb_seqr.sv"
`include "ahb_drv.sv"
`include "ahb_mon.sv"
`include "ahb_agt.sv"
`include "ahb_agt_top.sv"

`include "apb_config.sv"
`include "apb_trans.sv"
`include "apb_seqr.sv"
`include "apb_driver.sv"
`include "apb_mon.sv"
`include "apb_agt.sv"
`include "apb_agt_top.sv"

`include "env_config.sv"
`include "SB.sv"
`include "env.sv"
`include "test.sv"

endpackage
